`define DATA_WIDTH 32
`define ADDR_WIDTH 26
`define G_HISTORY_BITS 12

`define ROB_DEPTH 4
`define ROB_DEPTH_BITS 2

`define ALU_RES_STAT_DEPTH 4
`define ALU_RES_STAT_DEPTH_BITS 2

`define MEM_RES_STAT_DEPTH 4
`define MEM_RES_STAT_DEPTH_BITS 2

`define INSTRUCTION_QUEUE_DEPTH 4
`define INSTRUCTION_QUEUE_DEPTH_BITS 2

`define CHECKPOINT_BUFFER_DEPTH 4
`define CHECKPOINT_BUFFER_DEPTH_BITS 2


import mips_core_pkg::*;
