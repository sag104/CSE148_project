`define DATA_WIDTH 32
`define ADDR_WIDTH 26
`define G_HISTORY_BITS 12

import mips_core_pkg::*;
