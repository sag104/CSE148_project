import mips_core_pkg::*;
