`define DATA_WIDTH 32
`define ADDR_WIDTH 26

import mips_core_pkg::*;
