`define DATA_WIDTH 32
`define ADDR_WIDTH 26
`define G_HISTORY_BITS 12
`define ROB_DEPTH 4
`define RESERVATION_STATION_DEPTH 4

import mips_core_pkg::*;
